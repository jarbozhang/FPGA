// syncfifo_showahead_sclr_w8d64.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module syncfifo_showahead_sclr_w8d64 (
		input  wire [7:0] data,         //  fifo_input.datain
		input  wire       wrreq,        //            .wrreq
		input  wire       rdreq,        //            .rdreq
		input  wire       clock,        //            .clk
		input  wire       sclr,         //            .sclr
		output wire [7:0] q,            // fifo_output.dataout
		output wire [5:0] usedw,        //            .usedw
		output wire       full,         //            .full
		output wire       empty,        //            .empty
		output wire       almost_empty  //            .almost_empty
	);

	syncfifo_showahead_sclr_w8d64_fifo_191_qw52ykq fifo_0 (
		.data         (data),         //  fifo_input.datain
		.wrreq        (wrreq),        //            .wrreq
		.rdreq        (rdreq),        //            .rdreq
		.clock        (clock),        //            .clk
		.sclr         (sclr),         //            .sclr
		.q            (q),            // fifo_output.dataout
		.usedw        (usedw),        //            .usedw
		.full         (full),         //            .full
		.empty        (empty),        //            .empty
		.almost_empty (almost_empty)  //            .almost_empty
	);

endmodule
